// ALU to perform add, subtract, multiply and divide
module ALU(
    data1_i,
    data2_i,
    ALU_Ctrl_i,
    data_o,
    Zero_o
);

// Ports
// Wires and Registers

endmodule
