// Adder to compute the next PC
module Adder(
    data1_in,
    data2_in,
    data_o
);

// Ports
// Wires and Registers

endmodule
