// MUX three values of length 32 bits
module MUX32(
    data1_i,
    data2_i,
    data3_i,
    select_i,
    data_o
);