// Shift the immediate left 1 and pass it to Adder.v
module Shifter(
    data_i,
    data_o
);

// Ports
input   [31:0]  data_i;
output  [31:0]  data_o;

// Wires and Registers

// Assignment

endmodule
