// Control unit sending control signals
module Control(
    Op_i,
    Branch_o,
    MemRead_o,
    MemtoReg_o,
    ALUOp_o,
    MemWrite_o,
    ALUSrc_o,
    RegWrite_o
);

// Ports
// Wires and Registers
// Assignment

endmodule
