// Sign extend the immediate and pass it to Shifter.v
module Sign_Extend(
    data_i,
    data_o
);

// Ports
input   [31:0]  data_i;
output  [31:0]  data_o;

// Wires and Registers

endmodule
