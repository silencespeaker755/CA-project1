module ALU_Control
(
	func_i,
	ALUOp_i,
	ALUCtrl_o
);

// Ports

input  [3:0]		func_i;
input  [1:0]		ALIOp_i;
output [2:0]		ALUCtrl_o;


// Wires and Registers

// Assignment

endmodule