// MUX three values of length 32 bits
module MUX32(
    RS1data_EX_i,
    RS2data_EX_i,
    RDdata_WB_i,
    data3_i,
    select_i,
    data_o
);